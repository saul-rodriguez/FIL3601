* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : opamp1                                       *
* Netlisted  : Wed Sep  3 16:39:08 2025                     *
* PVS Version: 24.11-s045 Mon Jan 27 22:18:54 PST 2025      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(nel) nel ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pel) pel pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 MOSVC() mosvc p1trm(G) nwtrm(NW) bulk(SB)
*.DEVTMPLT 3 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 4 R(rpp1k1_3) rpp1k1_n p1trm(POS) p1trm(NEG) nwtrm(SUB)
*.DEVTMPLT 5 C(cmm5t) cmim capm(POS) m4trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MOSVC                                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MOSVC G NW SB
.ends MOSVC

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_756917543330                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_756917543330 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
R0 2 1 L=0.00012448 W=2e-06 $[rpp1k1_3] $SUB=3 $X=-2220 $Y=0 $dt=4
.ends rpp1k1_3_CDNS_756917543330

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nel_CDNS_756917543331                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nel_CDNS_756917543331 1 2 3 4
** N=4 EP=4 FDC=16
M0 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=2.4e-12 PD=5.54e-06 PS=1.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=790 $Y=0 $dt=0
M2 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=1580 $Y=0 $dt=0
M3 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=2370 $Y=0 $dt=0
M4 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=3160 $Y=0 $dt=0
M5 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=3950 $Y=0 $dt=0
M6 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=4740 $Y=0 $dt=0
M7 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=5530 $Y=0 $dt=0
M8 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=6320 $Y=0 $dt=0
M9 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=7110 $Y=0 $dt=0
M10 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=7900 $Y=0 $dt=0
M11 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=8690 $Y=0 $dt=0
M12 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=9480 $Y=0 $dt=0
M13 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=10270 $Y=0 $dt=0
M14 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=11060 $Y=0 $dt=0
M15 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=2.4e-12 AS=1.35e-12 PD=1.096e-05 PS=5.54e-06 $X=11850 $Y=0 $dt=0
.ends nel_CDNS_756917543331

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nel_CDNS_756917543332                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nel_CDNS_756917543332 1 2 3
** N=3 EP=3 FDC=8
M0 2 2 1 3 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=2.4e-12 PD=5.54e-06 PS=1.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 2 3 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=790 $Y=0 $dt=0
M2 2 2 1 3 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=1580 $Y=0 $dt=0
M3 1 2 2 3 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=2370 $Y=0 $dt=0
M4 2 2 1 3 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=3160 $Y=0 $dt=0
M5 1 2 2 3 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=3950 $Y=0 $dt=0
M6 2 2 1 3 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=4740 $Y=0 $dt=0
M7 1 2 2 3 nel L=2.5e-07 W=5e-06 AD=2.4e-12 AS=1.35e-12 PD=1.096e-05 PS=5.54e-06 $X=5530 $Y=0 $dt=0
.ends nel_CDNS_756917543332

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pel_CDNS_756917543334                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pel_CDNS_756917543334 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=8
M0 3 2 1 1 pel L=5e-07 W=2.5e-06 AD=6.75e-13 AS=1.2e-12 PD=3.04e-06 PS=5.96e-06 $X=0 $Y=0 $dt=1
M1 1 2 3 1 pel L=5e-07 W=2.5e-06 AD=6.75e-13 AS=6.75e-13 PD=3.04e-06 PS=3.04e-06 $X=1040 $Y=0 $dt=1
M2 3 2 1 1 pel L=5e-07 W=2.5e-06 AD=6.75e-13 AS=6.75e-13 PD=3.04e-06 PS=3.04e-06 $X=2080 $Y=0 $dt=1
M3 1 2 3 1 pel L=5e-07 W=2.5e-06 AD=6.75e-13 AS=6.75e-13 PD=3.04e-06 PS=3.04e-06 $X=3120 $Y=0 $dt=1
M4 3 2 1 1 pel L=5e-07 W=2.5e-06 AD=6.75e-13 AS=6.75e-13 PD=3.04e-06 PS=3.04e-06 $X=4160 $Y=0 $dt=1
M5 1 2 3 1 pel L=5e-07 W=2.5e-06 AD=6.75e-13 AS=6.75e-13 PD=3.04e-06 PS=3.04e-06 $X=5200 $Y=0 $dt=1
M6 3 2 1 1 pel L=5e-07 W=2.5e-06 AD=6.75e-13 AS=6.75e-13 PD=3.04e-06 PS=3.04e-06 $X=6240 $Y=0 $dt=1
M7 1 2 3 1 pel L=5e-07 W=2.5e-06 AD=1.2e-12 AS=6.75e-13 PD=5.96e-06 PS=3.04e-06 $X=7280 $Y=0 $dt=1
.ends pel_CDNS_756917543334

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nel_CDNS_756917543335                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nel_CDNS_756917543335 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 nel L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends nel_CDNS_756917543335

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pel_CDNS_756917543336                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pel_CDNS_756917543336 1 2 3
*.DEVICECLIMB
** N=4 EP=3 FDC=1
M0 3 2 1 1 pel L=2e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pel_CDNS_756917543336

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mosvc_CDNS_756917543339                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mosvc_CDNS_756917543339 1 2
** N=2 EP=2 FDC=2
X0 2 1 1 MOSVC w=8e-06 l=1e-05 $X=0 $Y=0 $dt=2
D1 1 1 p_dnw AREA=1.9232e-11 PJ=4.012e-05 perimeter=4.012e-05 $X=-600 $Y=-430 $dt=3
.ends mosvc_CDNS_756917543339

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mosvc_CDNS_7569175433310                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mosvc_CDNS_7569175433310 1 2
** N=2 EP=2 FDC=2
X0 2 1 1 MOSVC w=1.8e-05 l=1e-05 $X=0 $Y=0 $dt=2
D1 1 1 p_dnw AREA=3.1232e-11 PJ=6.012e-05 perimeter=6.012e-05 $X=-600 $Y=-430 $dt=3
.ends mosvc_CDNS_7569175433310

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nel_CDNS_756917543338                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nel_CDNS_756917543338 1
** N=1 EP=1 FDC=1
M0 1 1 1 1 nel L=2e-06 W=1e-06 AD=4.8e-13 AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 $X=0 $Y=0 $dt=0
.ends nel_CDNS_756917543338

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A1 1
** N=1 EP=1 FDC=2
X0 1 nel_CDNS_756917543338 $T=740 350 0 0 $X=0 $Y=0
X1 1 nel_CDNS_756917543338 $T=3980 350 0 0 $X=3240 $Y=0
.ends MASCO__A1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nel_CDNS_756917543337                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nel_CDNS_756917543337 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 nel L=2e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends nel_CDNS_756917543337

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A2 1 2 3 4 5
** N=5 EP=5 FDC=2
X0 1 2 3 nel_CDNS_756917543337 $T=740 350 0 0 $X=0 $Y=0
X1 1 4 5 nel_CDNS_756917543337 $T=3980 350 0 0 $X=3240 $Y=0
.ends MASCO__A2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A3                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A3 1 2 3 4 5 6
** N=6 EP=6 FDC=4
X0 1 2 3 4 5 MASCO__A2 $T=0 0 0 0 $X=0 $Y=0
X1 1 4 6 4 6 MASCO__A2 $T=6480 0 0 0 $X=6480 $Y=0
.ends MASCO__A3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: opamp1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt opamp1 BIAS GNDA INN INP OUT VDDA
** N=12 EP=6 FDC=156
X391 2 12 VDDA rpp1k1_3_CDNS_756917543330 $T=71840 92685 1 270 $X=49280 $Y=80495
X392 7 BIAS 4 GNDA nel_CDNS_756917543331 $T=31115 23480 1 0 $X=30375 $Y=17910
X393 5 BIAS GNDA nel_CDNS_756917543332 $T=18470 23480 1 0 $X=17730 $Y=17910
X394 VDDA 2 OUT pel_CDNS_756917543334 $T=57470 103255 0 180 $X=48780 $Y=100185
X395 GNDA GNDA GNDA GNDA nel_CDNS_756917543335 $T=12080 38620 0 0 $X=11340 $Y=38270
X396 GNDA GNDA GNDA GNDA nel_CDNS_756917543335 $T=12080 61580 1 0 $X=11340 $Y=51010
X397 4 INN 3 GNDA nel_CDNS_756917543335 $T=14320 38620 0 0 $X=13580 $Y=38270
X398 4 INP 2 GNDA nel_CDNS_756917543335 $T=14320 61580 1 0 $X=13580 $Y=51010
X399 4 INP 2 GNDA nel_CDNS_756917543335 $T=16560 38620 0 0 $X=15820 $Y=38270
X400 4 INN 3 GNDA nel_CDNS_756917543335 $T=16560 61580 1 0 $X=15820 $Y=51010
X401 4 INN 3 GNDA nel_CDNS_756917543335 $T=18800 38620 0 0 $X=18060 $Y=38270
X402 4 INP 2 GNDA nel_CDNS_756917543335 $T=18800 61580 1 0 $X=18060 $Y=51010
X403 4 INP 2 GNDA nel_CDNS_756917543335 $T=21040 38620 0 0 $X=20300 $Y=38270
X404 4 INN 3 GNDA nel_CDNS_756917543335 $T=21040 61580 1 0 $X=20300 $Y=51010
X405 4 INN 3 GNDA nel_CDNS_756917543335 $T=23280 38620 0 0 $X=22540 $Y=38270
X406 4 INP 2 GNDA nel_CDNS_756917543335 $T=23280 61580 1 0 $X=22540 $Y=51010
X407 4 INP 2 GNDA nel_CDNS_756917543335 $T=25520 38620 0 0 $X=24780 $Y=38270
X408 4 INN 3 GNDA nel_CDNS_756917543335 $T=25520 61580 1 0 $X=24780 $Y=51010
X409 4 INN 3 GNDA nel_CDNS_756917543335 $T=27760 38620 0 0 $X=27020 $Y=38270
X410 4 INP 2 GNDA nel_CDNS_756917543335 $T=27760 61580 1 0 $X=27020 $Y=51010
X411 4 INP 2 GNDA nel_CDNS_756917543335 $T=30000 38620 0 0 $X=29260 $Y=38270
X412 4 INN 3 GNDA nel_CDNS_756917543335 $T=30000 61580 1 0 $X=29260 $Y=51010
X413 4 INN 3 GNDA nel_CDNS_756917543335 $T=32240 38620 0 0 $X=31500 $Y=38270
X414 4 INP 2 GNDA nel_CDNS_756917543335 $T=32240 61580 1 0 $X=31500 $Y=51010
X415 4 INP 2 GNDA nel_CDNS_756917543335 $T=34480 38620 0 0 $X=33740 $Y=38270
X416 4 INN 3 GNDA nel_CDNS_756917543335 $T=34480 61580 1 0 $X=33740 $Y=51010
X417 GNDA GNDA GNDA GNDA nel_CDNS_756917543335 $T=36720 38620 0 0 $X=35980 $Y=38270
X418 GNDA GNDA GNDA GNDA nel_CDNS_756917543335 $T=36720 61580 1 0 $X=35980 $Y=51010
X419 VDDA VDDA VDDA pel_CDNS_756917543336 $T=8410 79155 0 0 $X=7500 $Y=78725
X420 VDDA VDDA VDDA pel_CDNS_756917543336 $T=8410 101415 1 0 $X=7500 $Y=90845
X421 VDDA 3 2 pel_CDNS_756917543336 $T=11650 79155 0 0 $X=10740 $Y=78725
X422 VDDA 3 3 pel_CDNS_756917543336 $T=11650 101415 1 0 $X=10740 $Y=90845
X423 VDDA 3 3 pel_CDNS_756917543336 $T=14890 79155 0 0 $X=13980 $Y=78725
X424 VDDA 3 2 pel_CDNS_756917543336 $T=14890 101415 1 0 $X=13980 $Y=90845
X425 VDDA 3 2 pel_CDNS_756917543336 $T=18130 79155 0 0 $X=17220 $Y=78725
X426 VDDA 3 3 pel_CDNS_756917543336 $T=18130 101415 1 0 $X=17220 $Y=90845
X427 VDDA 3 3 pel_CDNS_756917543336 $T=21370 79155 0 0 $X=20460 $Y=78725
X428 VDDA 3 2 pel_CDNS_756917543336 $T=21370 101415 1 0 $X=20460 $Y=90845
X429 VDDA 3 3 pel_CDNS_756917543336 $T=24610 79155 0 0 $X=23700 $Y=78725
X430 VDDA 3 2 pel_CDNS_756917543336 $T=24610 101415 1 0 $X=23700 $Y=90845
X431 VDDA 3 2 pel_CDNS_756917543336 $T=27850 79155 0 0 $X=26940 $Y=78725
X432 VDDA 3 3 pel_CDNS_756917543336 $T=27850 101415 1 0 $X=26940 $Y=90845
X433 VDDA 3 3 pel_CDNS_756917543336 $T=31090 79155 0 0 $X=30180 $Y=78725
X434 VDDA 3 2 pel_CDNS_756917543336 $T=31090 101415 1 0 $X=30180 $Y=90845
X435 VDDA 3 2 pel_CDNS_756917543336 $T=34330 79155 0 0 $X=33420 $Y=78725
X436 VDDA 3 3 pel_CDNS_756917543336 $T=34330 101415 1 0 $X=33420 $Y=90845
X437 VDDA VDDA VDDA pel_CDNS_756917543336 $T=37570 79155 0 0 $X=36660 $Y=78725
X438 VDDA VDDA VDDA pel_CDNS_756917543336 $T=37570 101415 1 0 $X=36660 $Y=90845
X439 GNDA VDDA mosvc_CDNS_756917543339 $T=63350 99890 0 0 $X=62610 $Y=99460
X440 GNDA BIAS mosvc_CDNS_7569175433310 $T=2695 11965 0 0 $X=1955 $Y=11535
X441 GNDA MASCO__A1 $T=55180 17760 0 0 $X=55180 $Y=17760
X442 GNDA MASCO__A1 $T=55180 73640 0 0 $X=55180 $Y=73640
X443 GNDA MASCO__A1 $T=61660 17760 0 0 $X=61660 $Y=17760
X444 GNDA MASCO__A1 $T=61660 73640 0 0 $X=61660 $Y=73640
X445 GNDA MASCO__A1 $T=68140 17760 0 0 $X=68140 $Y=17760
X446 GNDA MASCO__A1 $T=68140 73640 0 0 $X=68140 $Y=73640
X447 GNDA MASCO__A1 $T=74620 17760 0 0 $X=74620 $Y=17760
X448 GNDA MASCO__A1 $T=74620 73640 0 0 $X=74620 $Y=73640
X449 GNDA MASCO__A1 $T=81100 17760 0 0 $X=81100 $Y=17760
X450 GNDA MASCO__A1 $T=81100 73640 0 0 $X=81100 $Y=73640
X451 GNDA MASCO__A1 $T=87580 17760 0 0 $X=87580 $Y=17760
X452 GNDA MASCO__A1 $T=87580 73640 0 0 $X=87580 $Y=73640
X453 GNDA MASCO__A1 $T=94060 17760 0 0 $X=94060 $Y=17760
X454 GNDA MASCO__A1 $T=94060 73640 0 0 $X=94060 $Y=73640
X455 GNDA 5 OUT GNDA GNDA MASCO__A2 $T=94060 24980 0 0 $X=94060 $Y=24980
X456 GNDA 5 OUT GNDA GNDA MASCO__A2 $T=94060 41200 0 0 $X=94060 $Y=41200
X457 GNDA 5 OUT GNDA GNDA MASCO__A2 $T=94060 57420 0 0 $X=94060 $Y=57420
X458 GNDA GNDA GNDA 5 OUT OUT MASCO__A3 $T=55180 24980 0 0 $X=55180 $Y=24980
X459 GNDA GNDA GNDA 5 OUT OUT MASCO__A3 $T=55180 41200 0 0 $X=55180 $Y=41200
X460 GNDA GNDA GNDA 5 OUT OUT MASCO__A3 $T=55180 57420 0 0 $X=55180 $Y=57420
X461 GNDA 5 OUT 5 OUT 7 MASCO__A3 $T=68140 24980 0 0 $X=68140 $Y=24980
X462 GNDA 5 OUT 5 OUT 5 MASCO__A3 $T=68140 41200 0 0 $X=68140 $Y=41200
X463 GNDA 5 OUT 5 OUT 7 MASCO__A3 $T=68140 57420 0 0 $X=68140 $Y=57420
X464 GNDA 5 OUT 5 OUT OUT MASCO__A3 $T=81100 24980 0 0 $X=81100 $Y=24980
X465 GNDA 5 OUT 5 OUT OUT MASCO__A3 $T=81100 41200 0 0 $X=81100 $Y=41200
X466 GNDA 5 OUT 5 OUT OUT MASCO__A3 $T=81100 57420 0 0 $X=81100 $Y=57420
D0 GNDA VDDA p_dnw AREA=1.63313e-09 PJ=0.00016212 perimeter=0.00016212 $X=2180 $Y=71565 $dt=3
D1 GNDA VDDA p_dnw AREA=1.34725e-10 PJ=4.668e-05 perimeter=4.668e-05 $X=47140 $Y=98545 $dt=3
D2 GNDA VDDA p_dnw AREA=4.85498e-10 PJ=8.938e-05 perimeter=8.938e-05 $X=47640 $Y=78855 $dt=3
D3 GNDA VDDA p_dnw AREA=1.00372e-09 PJ=0.00012712 perimeter=0.00012712 $X=75350 $Y=79725 $dt=3
C4 12 OUT area=7.5e-10 perimeter=0.00011 $[cmm5t] $X=77490 $Y=81865 $dt=5
.ends opamp1
