* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* CDL Netlist:                                              *
*                                                           *
* Cell Name  : opamp1                                       *
* Netlisted  : Wed Sep  3 16:39:08 2025                     *
* PVS Version: 24.11-s045 Mon Jan 27 22:18:54 PST 2025      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
*.LDD
*.DEVTMPLT 0 MN(nel) nel ndiff(D) p1trm(G) ndiff(S) bulk(B)
*.DEVTMPLT 1 MP(pel) pel pdiff(D) p1trm(G) pdiff(S) nwtrm(B)
*.DEVTMPLT 2 MOSVC() mosvc p1trm(G) nwtrm(NW) bulk(SB)
*.DEVTMPLT 3 D(p_dnw) p_dnw bulk(POS) nwtrm(NEG)
*.DEVTMPLT 4 R(rpp1k1_3) rpp1k1_n p1trm(POS) p1trm(NEG) nwtrm(SUB)
*.DEVTMPLT 5 C(cmm5t) cmim capm(POS) m4trm(NEG)

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_756917543330                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_756917543330 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_756917543330

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_756917543331                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_756917543331 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_756917543331

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_756917543332                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_756917543332 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_756917543332

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_756917543334                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_756917543334 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_756917543334

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_756917543336                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_756917543336 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_756917543336

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_756917543338                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_756917543338 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_756917543338

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA1_C_CDNS_756917543339                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA1_C_CDNS_756917543339 1
** N=1 EP=1 FDC=0
.ends VIA1_C_CDNS_756917543339

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: VIA2_C_CDNS_7569175433317                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt VIA2_C_CDNS_7569175433317 1
** N=1 EP=1 FDC=0
.ends VIA2_C_CDNS_7569175433317

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: rpp1k1_3_CDNS_756917543330                      *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt rpp1k1_3_CDNS_756917543330 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
R0 2 1 L=0.00012448 W=2e-06 $[rpp1k1_3] $SUB=3 $X=-2220 $Y=0 $dt=4
.ends rpp1k1_3_CDNS_756917543330

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nel_CDNS_756917543331                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nel_CDNS_756917543331 1 2 3 4
** N=4 EP=4 FDC=16
M0 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=2.4e-12 PD=5.54e-06 PS=1.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=790 $Y=0 $dt=0
M2 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=1580 $Y=0 $dt=0
M3 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=2370 $Y=0 $dt=0
M4 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=3160 $Y=0 $dt=0
M5 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=3950 $Y=0 $dt=0
M6 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=4740 $Y=0 $dt=0
M7 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=5530 $Y=0 $dt=0
M8 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=6320 $Y=0 $dt=0
M9 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=7110 $Y=0 $dt=0
M10 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=7900 $Y=0 $dt=0
M11 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=8690 $Y=0 $dt=0
M12 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=9480 $Y=0 $dt=0
M13 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=10270 $Y=0 $dt=0
M14 3 2 1 4 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=11060 $Y=0 $dt=0
M15 1 2 3 4 nel L=2.5e-07 W=5e-06 AD=2.4e-12 AS=1.35e-12 PD=1.096e-05 PS=5.54e-06 $X=11850 $Y=0 $dt=0
.ends nel_CDNS_756917543331

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nel_CDNS_756917543332                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nel_CDNS_756917543332 1 2 3
** N=3 EP=3 FDC=8
M0 2 2 1 3 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=2.4e-12 PD=5.54e-06 PS=1.096e-05 $X=0 $Y=0 $dt=0
M1 1 2 2 3 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=790 $Y=0 $dt=0
M2 2 2 1 3 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=1580 $Y=0 $dt=0
M3 1 2 2 3 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=2370 $Y=0 $dt=0
M4 2 2 1 3 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=3160 $Y=0 $dt=0
M5 1 2 2 3 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=3950 $Y=0 $dt=0
M6 2 2 1 3 nel L=2.5e-07 W=5e-06 AD=1.35e-12 AS=1.35e-12 PD=5.54e-06 PS=5.54e-06 $X=4740 $Y=0 $dt=0
M7 1 2 2 3 nel L=2.5e-07 W=5e-06 AD=2.4e-12 AS=1.35e-12 PD=1.096e-05 PS=5.54e-06 $X=5530 $Y=0 $dt=0
.ends nel_CDNS_756917543332

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pel_CDNS_756917543334                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pel_CDNS_756917543334 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=8
M0 3 2 1 1 pel L=5e-07 W=2.5e-06 AD=6.75e-13 AS=1.2e-12 PD=3.04e-06 PS=5.96e-06 $X=0 $Y=0 $dt=1
M1 1 2 3 1 pel L=5e-07 W=2.5e-06 AD=6.75e-13 AS=6.75e-13 PD=3.04e-06 PS=3.04e-06 $X=1040 $Y=0 $dt=1
M2 3 2 1 1 pel L=5e-07 W=2.5e-06 AD=6.75e-13 AS=6.75e-13 PD=3.04e-06 PS=3.04e-06 $X=2080 $Y=0 $dt=1
M3 1 2 3 1 pel L=5e-07 W=2.5e-06 AD=6.75e-13 AS=6.75e-13 PD=3.04e-06 PS=3.04e-06 $X=3120 $Y=0 $dt=1
M4 3 2 1 1 pel L=5e-07 W=2.5e-06 AD=6.75e-13 AS=6.75e-13 PD=3.04e-06 PS=3.04e-06 $X=4160 $Y=0 $dt=1
M5 1 2 3 1 pel L=5e-07 W=2.5e-06 AD=6.75e-13 AS=6.75e-13 PD=3.04e-06 PS=3.04e-06 $X=5200 $Y=0 $dt=1
M6 3 2 1 1 pel L=5e-07 W=2.5e-06 AD=6.75e-13 AS=6.75e-13 PD=3.04e-06 PS=3.04e-06 $X=6240 $Y=0 $dt=1
M7 1 2 3 1 pel L=5e-07 W=2.5e-06 AD=1.2e-12 AS=6.75e-13 PD=5.96e-06 PS=3.04e-06 $X=7280 $Y=0 $dt=1
.ends pel_CDNS_756917543334

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nel_CDNS_756917543335                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nel_CDNS_756917543335 1 2 3 4
** N=4 EP=4 FDC=1
M0 3 2 1 4 nel L=1e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends nel_CDNS_756917543335

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: pel_CDNS_756917543336                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt pel_CDNS_756917543336 1 2 3 4
*.DEVICECLIMB
** N=4 EP=4 FDC=1
M0 3 2 1 1 pel L=2e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=1
.ends pel_CDNS_756917543336

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mosvc_CDNS_756917543339                         *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mosvc_CDNS_756917543339 1 2
** N=2 EP=2 FDC=2
X0 2 1 1 MOSVC w=8e-06 l=1e-05 $X=0 $Y=0 $dt=2
D1 1 1 p_dnw AREA=1.9232e-11 PJ=4.012e-05 perimeter=4.012e-05 $X=-600 $Y=-430 $dt=3
.ends mosvc_CDNS_756917543339

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: mosvc_CDNS_7569175433310                        *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt mosvc_CDNS_7569175433310 1 2
** N=2 EP=2 FDC=2
X0 2 1 1 MOSVC w=1.8e-05 l=1e-05 $X=0 $Y=0 $dt=2
D1 1 1 p_dnw AREA=3.1232e-11 PJ=6.012e-05 perimeter=6.012e-05 $X=-600 $Y=-430 $dt=3
.ends mosvc_CDNS_7569175433310

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nel_CDNS_756917543338                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nel_CDNS_756917543338 1
** N=1 EP=1 FDC=1
M0 1 1 1 1 nel L=2e-06 W=1e-06 AD=4.8e-13 AS=4.8e-13 PD=2.96e-06 PS=2.96e-06 $X=0 $Y=0 $dt=0
.ends nel_CDNS_756917543338

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A1                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A1 1
** N=1 EP=1 FDC=2
X0 1 nel_CDNS_756917543338 $T=740 350 0 0 $X=0 $Y=0
X1 1 nel_CDNS_756917543338 $T=3980 350 0 0 $X=3240 $Y=0
.ends MASCO__A1

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: nel_CDNS_756917543337                           *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt nel_CDNS_756917543337 1 2 3
** N=3 EP=3 FDC=1
M0 3 2 1 1 nel L=2e-06 W=1e-05 AD=4.8e-12 AS=4.8e-12 PD=2.096e-05 PS=2.096e-05 $X=0 $Y=0 $dt=0
.ends nel_CDNS_756917543337

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A2                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A2 1 2 3 4 5
** N=5 EP=5 FDC=2
X0 1 2 3 nel_CDNS_756917543337 $T=740 350 0 0 $X=0 $Y=0
X1 1 4 5 nel_CDNS_756917543337 $T=3980 350 0 0 $X=3240 $Y=0
.ends MASCO__A2

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: MASCO__A3                                       *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt MASCO__A3 1 2 3 4 5 6
** N=6 EP=6 FDC=4
X0 1 2 3 4 5 MASCO__A2 $T=0 0 0 0 $X=0 $Y=0
X1 1 4 6 4 6 MASCO__A2 $T=6480 0 0 0 $X=6480 $Y=0
.ends MASCO__A3

* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
* Sub cell: opamp1                                          *
* +++++++++++++++++++++++++++++++++++++++++++++++++++++++++ *
.subckt opamp1 6 11 9 10 8 1
** N=12 EP=6 FDC=156
X0 1 VIA1_C_CDNS_756917543330 $T=8140 77635 0 0 $X=8000 $Y=76925
X1 1 VIA1_C_CDNS_756917543330 $T=8140 102935 0 0 $X=8000 $Y=102225
X2 1 VIA1_C_CDNS_756917543330 $T=10680 77635 0 0 $X=10540 $Y=76925
X3 1 VIA1_C_CDNS_756917543330 $T=10680 102935 0 0 $X=10540 $Y=102225
X4 1 VIA1_C_CDNS_756917543330 $T=11380 77635 0 0 $X=11240 $Y=76925
X5 1 VIA1_C_CDNS_756917543330 $T=11380 102935 0 0 $X=11240 $Y=102225
X6 2 VIA1_C_CDNS_756917543330 $T=13920 75795 0 0 $X=13780 $Y=75085
X7 3 VIA1_C_CDNS_756917543330 $T=13920 104775 0 0 $X=13780 $Y=104065
X8 4 VIA1_C_CDNS_756917543330 $T=14050 37180 0 0 $X=13910 $Y=36470
X9 4 VIA1_C_CDNS_756917543330 $T=14050 63020 0 0 $X=13910 $Y=62310
X10 1 VIA1_C_CDNS_756917543330 $T=14620 77635 0 0 $X=14480 $Y=76925
X11 1 VIA1_C_CDNS_756917543330 $T=14620 102935 0 0 $X=14480 $Y=102225
X12 3 VIA1_C_CDNS_756917543330 $T=15590 35340 0 0 $X=15450 $Y=34630
X13 2 VIA1_C_CDNS_756917543330 $T=15590 64860 0 0 $X=15450 $Y=64150
X14 4 VIA1_C_CDNS_756917543330 $T=16290 37180 0 0 $X=16150 $Y=36470
X15 4 VIA1_C_CDNS_756917543330 $T=16290 63020 0 0 $X=16150 $Y=62310
X16 3 VIA1_C_CDNS_756917543330 $T=17160 73955 0 0 $X=17020 $Y=73245
X17 2 VIA1_C_CDNS_756917543330 $T=17160 106615 0 0 $X=17020 $Y=105905
X18 2 VIA1_C_CDNS_756917543330 $T=17830 33500 0 0 $X=17690 $Y=32790
X19 3 VIA1_C_CDNS_756917543330 $T=17830 66700 0 0 $X=17690 $Y=65990
X20 1 VIA1_C_CDNS_756917543330 $T=17860 77635 0 0 $X=17720 $Y=76925
X21 1 VIA1_C_CDNS_756917543330 $T=17860 102935 0 0 $X=17720 $Y=102225
X22 5 VIA1_C_CDNS_756917543330 $T=18200 24920 1 0 $X=18060 $Y=24210
X23 4 VIA1_C_CDNS_756917543330 $T=18530 37180 0 0 $X=18390 $Y=36470
X24 4 VIA1_C_CDNS_756917543330 $T=18530 63020 0 0 $X=18390 $Y=62310
X25 6 VIA1_C_CDNS_756917543330 $T=18990 26760 1 0 $X=18850 $Y=26050
X26 5 VIA1_C_CDNS_756917543330 $T=19780 24920 1 0 $X=19640 $Y=24210
X27 3 VIA1_C_CDNS_756917543330 $T=20070 35340 0 0 $X=19930 $Y=34630
X28 2 VIA1_C_CDNS_756917543330 $T=20070 64860 0 0 $X=19930 $Y=64150
X29 2 VIA1_C_CDNS_756917543330 $T=20400 75795 0 0 $X=20260 $Y=75085
X30 3 VIA1_C_CDNS_756917543330 $T=20400 104775 0 0 $X=20260 $Y=104065
X31 6 VIA1_C_CDNS_756917543330 $T=20570 26760 1 0 $X=20430 $Y=26050
X32 4 VIA1_C_CDNS_756917543330 $T=20770 37180 0 0 $X=20630 $Y=36470
X33 4 VIA1_C_CDNS_756917543330 $T=20770 63020 0 0 $X=20630 $Y=62310
X34 1 VIA1_C_CDNS_756917543330 $T=21100 77635 0 0 $X=20960 $Y=76925
X35 1 VIA1_C_CDNS_756917543330 $T=21100 102935 0 0 $X=20960 $Y=102225
X36 5 VIA1_C_CDNS_756917543330 $T=21360 24920 1 0 $X=21220 $Y=24210
X37 6 VIA1_C_CDNS_756917543330 $T=22150 26760 1 0 $X=22010 $Y=26050
X38 2 VIA1_C_CDNS_756917543330 $T=22310 33500 0 0 $X=22170 $Y=32790
X39 3 VIA1_C_CDNS_756917543330 $T=22310 66700 0 0 $X=22170 $Y=65990
X40 5 VIA1_C_CDNS_756917543330 $T=22940 24920 1 0 $X=22800 $Y=24210
X41 4 VIA1_C_CDNS_756917543330 $T=23010 37180 0 0 $X=22870 $Y=36470
X42 4 VIA1_C_CDNS_756917543330 $T=23010 63020 0 0 $X=22870 $Y=62310
X43 3 VIA1_C_CDNS_756917543330 $T=23640 73955 0 0 $X=23500 $Y=73245
X44 2 VIA1_C_CDNS_756917543330 $T=23640 106615 0 0 $X=23500 $Y=105905
X45 6 VIA1_C_CDNS_756917543330 $T=23730 26760 1 0 $X=23590 $Y=26050
X46 1 VIA1_C_CDNS_756917543330 $T=24340 77635 0 0 $X=24200 $Y=76925
X47 1 VIA1_C_CDNS_756917543330 $T=24340 102935 0 0 $X=24200 $Y=102225
X48 5 VIA1_C_CDNS_756917543330 $T=24520 24920 1 0 $X=24380 $Y=24210
X49 3 VIA1_C_CDNS_756917543330 $T=24550 35340 0 0 $X=24410 $Y=34630
X50 2 VIA1_C_CDNS_756917543330 $T=24550 64860 0 0 $X=24410 $Y=64150
X51 4 VIA1_C_CDNS_756917543330 $T=25250 37180 0 0 $X=25110 $Y=36470
X52 4 VIA1_C_CDNS_756917543330 $T=25250 63020 0 0 $X=25110 $Y=62310
X53 2 VIA1_C_CDNS_756917543330 $T=26790 33500 0 0 $X=26650 $Y=32790
X54 3 VIA1_C_CDNS_756917543330 $T=26790 66700 0 0 $X=26650 $Y=65990
X55 3 VIA1_C_CDNS_756917543330 $T=26880 73955 0 0 $X=26740 $Y=73245
X56 2 VIA1_C_CDNS_756917543330 $T=26880 106615 0 0 $X=26740 $Y=105905
X57 4 VIA1_C_CDNS_756917543330 $T=27490 37180 0 0 $X=27350 $Y=36470
X58 4 VIA1_C_CDNS_756917543330 $T=27490 63020 0 0 $X=27350 $Y=62310
X59 1 VIA1_C_CDNS_756917543330 $T=27580 77635 0 0 $X=27440 $Y=76925
X60 1 VIA1_C_CDNS_756917543330 $T=27580 102935 0 0 $X=27440 $Y=102225
X61 3 VIA1_C_CDNS_756917543330 $T=29030 35340 0 0 $X=28890 $Y=34630
X62 2 VIA1_C_CDNS_756917543330 $T=29030 64860 0 0 $X=28890 $Y=64150
X63 4 VIA1_C_CDNS_756917543330 $T=29730 37180 0 0 $X=29590 $Y=36470
X64 4 VIA1_C_CDNS_756917543330 $T=29730 63020 0 0 $X=29590 $Y=62310
X65 2 VIA1_C_CDNS_756917543330 $T=30120 75795 0 0 $X=29980 $Y=75085
X66 3 VIA1_C_CDNS_756917543330 $T=30120 104775 0 0 $X=29980 $Y=104065
X67 1 VIA1_C_CDNS_756917543330 $T=30820 77635 0 0 $X=30680 $Y=76925
X68 1 VIA1_C_CDNS_756917543330 $T=30820 102935 0 0 $X=30680 $Y=102225
X69 7 VIA1_C_CDNS_756917543330 $T=30845 24920 1 0 $X=30705 $Y=24210
X70 2 VIA1_C_CDNS_756917543330 $T=31270 33500 0 0 $X=31130 $Y=32790
X71 3 VIA1_C_CDNS_756917543330 $T=31270 66700 0 0 $X=31130 $Y=65990
X72 4 VIA1_C_CDNS_756917543330 $T=31635 26760 1 0 $X=31495 $Y=26050
X73 4 VIA1_C_CDNS_756917543330 $T=31970 37180 0 0 $X=31830 $Y=36470
X74 4 VIA1_C_CDNS_756917543330 $T=31970 63020 0 0 $X=31830 $Y=62310
X75 7 VIA1_C_CDNS_756917543330 $T=32425 24920 1 0 $X=32285 $Y=24210
X76 4 VIA1_C_CDNS_756917543330 $T=33215 26760 1 0 $X=33075 $Y=26050
X77 3 VIA1_C_CDNS_756917543330 $T=33360 73955 0 0 $X=33220 $Y=73245
X78 2 VIA1_C_CDNS_756917543330 $T=33360 106615 0 0 $X=33220 $Y=105905
X79 3 VIA1_C_CDNS_756917543330 $T=33510 35340 0 0 $X=33370 $Y=34630
X80 2 VIA1_C_CDNS_756917543330 $T=33510 64860 0 0 $X=33370 $Y=64150
X81 7 VIA1_C_CDNS_756917543330 $T=34005 24920 1 0 $X=33865 $Y=24210
X82 1 VIA1_C_CDNS_756917543330 $T=34060 77635 0 0 $X=33920 $Y=76925
X83 1 VIA1_C_CDNS_756917543330 $T=34060 102935 0 0 $X=33920 $Y=102225
X84 4 VIA1_C_CDNS_756917543330 $T=34210 37180 0 0 $X=34070 $Y=36470
X85 4 VIA1_C_CDNS_756917543330 $T=34210 63020 0 0 $X=34070 $Y=62310
X86 4 VIA1_C_CDNS_756917543330 $T=34795 26760 1 0 $X=34655 $Y=26050
X87 7 VIA1_C_CDNS_756917543330 $T=35585 24920 1 0 $X=35445 $Y=24210
X88 2 VIA1_C_CDNS_756917543330 $T=35750 33500 0 0 $X=35610 $Y=32790
X89 3 VIA1_C_CDNS_756917543330 $T=35750 66700 0 0 $X=35610 $Y=65990
X90 4 VIA1_C_CDNS_756917543330 $T=36375 26760 1 0 $X=36235 $Y=26050
X91 2 VIA1_C_CDNS_756917543330 $T=36600 75795 0 0 $X=36460 $Y=75085
X92 3 VIA1_C_CDNS_756917543330 $T=36600 104775 0 0 $X=36460 $Y=104065
X93 7 VIA1_C_CDNS_756917543330 $T=37165 24920 1 0 $X=37025 $Y=24210
X94 1 VIA1_C_CDNS_756917543330 $T=37300 77635 0 0 $X=37160 $Y=76925
X95 1 VIA1_C_CDNS_756917543330 $T=37300 102935 0 0 $X=37160 $Y=102225
X96 4 VIA1_C_CDNS_756917543330 $T=37955 26760 1 0 $X=37815 $Y=26050
X97 7 VIA1_C_CDNS_756917543330 $T=38745 24920 1 0 $X=38605 $Y=24210
X98 4 VIA1_C_CDNS_756917543330 $T=39535 26760 1 0 $X=39395 $Y=26050
X99 1 VIA1_C_CDNS_756917543330 $T=39840 77635 0 0 $X=39700 $Y=76925
X100 1 VIA1_C_CDNS_756917543330 $T=39840 102935 0 0 $X=39700 $Y=102225
X101 7 VIA1_C_CDNS_756917543330 $T=40325 24920 1 0 $X=40185 $Y=24210
X102 4 VIA1_C_CDNS_756917543330 $T=41115 26760 1 0 $X=40975 $Y=26050
X103 7 VIA1_C_CDNS_756917543330 $T=41905 24920 1 0 $X=41765 $Y=24210
X104 4 VIA1_C_CDNS_756917543330 $T=42695 26760 1 0 $X=42555 $Y=26050
X105 7 VIA1_C_CDNS_756917543330 $T=43485 24920 1 0 $X=43345 $Y=24210
X106 1 VIA1_C_CDNS_756917543330 $T=49420 104775 0 180 $X=49280 $Y=104065
X107 8 VIA1_C_CDNS_756917543330 $T=50460 106615 0 180 $X=50320 $Y=105905
X108 1 VIA1_C_CDNS_756917543330 $T=51500 104775 0 180 $X=51360 $Y=104065
X109 8 VIA1_C_CDNS_756917543330 $T=52540 106615 0 180 $X=52400 $Y=105905
X110 1 VIA1_C_CDNS_756917543330 $T=53580 104775 0 180 $X=53440 $Y=104065
X111 8 VIA1_C_CDNS_756917543330 $T=54620 106615 0 180 $X=54480 $Y=105905
X112 1 VIA1_C_CDNS_756917543330 $T=55660 104775 0 180 $X=55520 $Y=104065
X113 8 VIA1_C_CDNS_756917543330 $T=56700 106615 0 180 $X=56560 $Y=105905
X114 1 VIA1_C_CDNS_756917543330 $T=57740 104775 0 180 $X=57600 $Y=104065
X115 2 VIA2_C_CDNS_756917543331 $T=4570 75795 0 0 $X=3860 $Y=75135
X116 2 VIA2_C_CDNS_756917543331 $T=4570 106615 0 0 $X=3860 $Y=105955
X117 1 VIA2_C_CDNS_756917543331 $T=6410 77635 0 0 $X=5700 $Y=76975
X118 1 VIA2_C_CDNS_756917543331 $T=6410 102935 0 0 $X=5700 $Y=102275
X119 2 VIA2_C_CDNS_756917543331 $T=6570 33500 0 0 $X=5860 $Y=32840
X120 2 VIA2_C_CDNS_756917543331 $T=6570 64860 0 0 $X=5860 $Y=64200
X121 3 VIA2_C_CDNS_756917543331 $T=8410 35340 0 0 $X=7700 $Y=34680
X122 3 VIA2_C_CDNS_756917543331 $T=8410 66700 0 0 $X=7700 $Y=66040
X123 4 VIA2_C_CDNS_756917543331 $T=10250 37180 0 0 $X=9540 $Y=36520
X124 4 VIA2_C_CDNS_756917543331 $T=10250 63020 0 0 $X=9540 $Y=62360
X125 4 VIA2_C_CDNS_756917543331 $T=39550 37180 0 0 $X=38840 $Y=36520
X126 4 VIA2_C_CDNS_756917543331 $T=39550 63020 0 0 $X=38840 $Y=62360
X127 2 VIA2_C_CDNS_756917543331 $T=41390 33500 0 0 $X=40680 $Y=32840
X128 2 VIA2_C_CDNS_756917543331 $T=41390 64860 0 0 $X=40680 $Y=64200
X129 1 VIA2_C_CDNS_756917543331 $T=41570 77635 0 0 $X=40860 $Y=76975
X130 1 VIA2_C_CDNS_756917543331 $T=41570 102935 0 0 $X=40860 $Y=102275
X131 3 VIA2_C_CDNS_756917543331 $T=43230 35340 0 0 $X=42520 $Y=34680
X132 3 VIA2_C_CDNS_756917543331 $T=43230 66700 0 0 $X=42520 $Y=66040
X133 3 VIA2_C_CDNS_756917543331 $T=43410 73955 0 0 $X=42700 $Y=73295
X134 3 VIA2_C_CDNS_756917543331 $T=43410 104775 0 0 $X=42700 $Y=104115
X135 3 VIA1_C_CDNS_756917543332 $T=12650 90265 0 0 $X=12510 $Y=90075
X136 9 VIA1_C_CDNS_756917543332 $T=14820 49730 0 0 $X=14680 $Y=49540
X137 10 VIA1_C_CDNS_756917543332 $T=14820 50470 0 0 $X=14680 $Y=50280
X138 3 VIA1_C_CDNS_756917543332 $T=15890 90265 0 0 $X=15750 $Y=90075
X139 9 VIA1_C_CDNS_756917543332 $T=16720 49730 0 0 $X=16580 $Y=49540
X140 10 VIA1_C_CDNS_756917543332 $T=17400 50470 0 0 $X=17260 $Y=50280
X141 3 VIA1_C_CDNS_756917543332 $T=19130 90265 0 0 $X=18990 $Y=90075
X142 9 VIA1_C_CDNS_756917543332 $T=19300 49730 0 0 $X=19160 $Y=49540
X143 10 VIA1_C_CDNS_756917543332 $T=19300 50470 0 0 $X=19160 $Y=50280
X144 9 VIA1_C_CDNS_756917543332 $T=21200 49730 0 0 $X=21060 $Y=49540
X145 10 VIA1_C_CDNS_756917543332 $T=21880 50470 0 0 $X=21740 $Y=50280
X146 3 VIA1_C_CDNS_756917543332 $T=22370 90265 0 0 $X=22230 $Y=90075
X147 9 VIA1_C_CDNS_756917543332 $T=23780 49730 0 0 $X=23640 $Y=49540
X148 10 VIA1_C_CDNS_756917543332 $T=23780 50470 0 0 $X=23640 $Y=50280
X149 3 VIA1_C_CDNS_756917543332 $T=25610 90265 0 0 $X=25470 $Y=90075
X150 9 VIA1_C_CDNS_756917543332 $T=25680 49730 0 0 $X=25540 $Y=49540
X151 10 VIA1_C_CDNS_756917543332 $T=26360 50470 0 0 $X=26220 $Y=50280
X152 9 VIA1_C_CDNS_756917543332 $T=28260 49730 0 0 $X=28120 $Y=49540
X153 10 VIA1_C_CDNS_756917543332 $T=28260 50470 0 0 $X=28120 $Y=50280
X154 3 VIA1_C_CDNS_756917543332 $T=28850 90265 0 0 $X=28710 $Y=90075
X155 9 VIA1_C_CDNS_756917543332 $T=30160 49730 0 0 $X=30020 $Y=49540
X156 10 VIA1_C_CDNS_756917543332 $T=30840 50470 0 0 $X=30700 $Y=50280
X157 3 VIA1_C_CDNS_756917543332 $T=32090 90265 0 0 $X=31950 $Y=90075
X158 9 VIA1_C_CDNS_756917543332 $T=32740 49730 0 0 $X=32600 $Y=49540
X159 10 VIA1_C_CDNS_756917543332 $T=32740 50470 0 0 $X=32600 $Y=50280
X160 9 VIA1_C_CDNS_756917543332 $T=34640 49730 0 0 $X=34500 $Y=49540
X161 10 VIA1_C_CDNS_756917543332 $T=35320 50470 0 0 $X=35180 $Y=50280
X162 3 VIA1_C_CDNS_756917543332 $T=35330 90265 0 0 $X=35190 $Y=90075
X163 11 VIA1_C_CDNS_756917543334 $T=55650 17120 0 0 $X=55510 $Y=16670
X164 11 VIA1_C_CDNS_756917543334 $T=55650 24340 0 0 $X=55510 $Y=23890
X165 11 VIA1_C_CDNS_756917543334 $T=55650 40560 0 0 $X=55510 $Y=40110
X166 11 VIA1_C_CDNS_756917543334 $T=55650 56780 0 0 $X=55510 $Y=56330
X167 11 VIA1_C_CDNS_756917543334 $T=55650 73000 0 0 $X=55510 $Y=72550
X168 11 VIA1_C_CDNS_756917543334 $T=56920 24340 0 0 $X=56780 $Y=23890
X169 11 VIA1_C_CDNS_756917543334 $T=56920 40560 0 0 $X=56780 $Y=40110
X170 11 VIA1_C_CDNS_756917543334 $T=56920 56780 0 0 $X=56780 $Y=56330
X171 11 VIA1_C_CDNS_756917543334 $T=56920 73000 0 0 $X=56780 $Y=72550
X172 11 VIA1_C_CDNS_756917543334 $T=58190 17120 0 0 $X=58050 $Y=16670
X173 11 VIA1_C_CDNS_756917543334 $T=58190 24340 0 0 $X=58050 $Y=23890
X174 11 VIA1_C_CDNS_756917543334 $T=58190 40560 0 0 $X=58050 $Y=40110
X175 11 VIA1_C_CDNS_756917543334 $T=58190 56780 0 0 $X=58050 $Y=56330
X176 11 VIA1_C_CDNS_756917543334 $T=58190 73000 0 0 $X=58050 $Y=72550
X177 11 VIA1_C_CDNS_756917543334 $T=58890 17120 0 0 $X=58750 $Y=16670
X178 11 VIA1_C_CDNS_756917543334 $T=58890 24340 0 0 $X=58750 $Y=23890
X179 11 VIA1_C_CDNS_756917543334 $T=58890 40560 0 0 $X=58750 $Y=40110
X180 11 VIA1_C_CDNS_756917543334 $T=58890 56780 0 0 $X=58750 $Y=56330
X181 11 VIA1_C_CDNS_756917543334 $T=58890 73000 0 0 $X=58750 $Y=72550
X182 11 VIA1_C_CDNS_756917543334 $T=60160 24340 0 0 $X=60020 $Y=23890
X183 5 VIA1_C_CDNS_756917543334 $T=60160 36540 0 0 $X=60020 $Y=36090
X184 5 VIA1_C_CDNS_756917543334 $T=60160 52760 0 0 $X=60020 $Y=52310
X185 5 VIA1_C_CDNS_756917543334 $T=60160 68980 0 0 $X=60020 $Y=68530
X186 11 VIA1_C_CDNS_756917543334 $T=61430 17120 0 0 $X=61290 $Y=16670
X187 8 VIA1_C_CDNS_756917543334 $T=61430 21660 0 0 $X=61290 $Y=21210
X188 8 VIA1_C_CDNS_756917543334 $T=61430 37880 0 0 $X=61290 $Y=37430
X189 8 VIA1_C_CDNS_756917543334 $T=61430 54100 0 0 $X=61290 $Y=53650
X190 11 VIA1_C_CDNS_756917543334 $T=61430 73000 0 0 $X=61290 $Y=72550
X191 11 VIA1_C_CDNS_756917543334 $T=62130 17120 0 0 $X=61990 $Y=16670
X192 11 VIA1_C_CDNS_756917543334 $T=62130 24340 0 0 $X=61990 $Y=23890
X193 11 VIA1_C_CDNS_756917543334 $T=62130 40560 0 0 $X=61990 $Y=40110
X194 11 VIA1_C_CDNS_756917543334 $T=62130 56780 0 0 $X=61990 $Y=56330
X195 11 VIA1_C_CDNS_756917543334 $T=62130 73000 0 0 $X=61990 $Y=72550
X196 11 VIA1_C_CDNS_756917543334 $T=63400 24340 0 0 $X=63260 $Y=23890
X197 5 VIA1_C_CDNS_756917543334 $T=63400 36540 0 0 $X=63260 $Y=36090
X198 5 VIA1_C_CDNS_756917543334 $T=63400 52760 0 0 $X=63260 $Y=52310
X199 5 VIA1_C_CDNS_756917543334 $T=63400 68980 0 0 $X=63260 $Y=68530
X200 11 VIA1_C_CDNS_756917543334 $T=64670 17120 0 0 $X=64530 $Y=16670
X201 8 VIA1_C_CDNS_756917543334 $T=64670 21660 0 0 $X=64530 $Y=21210
X202 8 VIA1_C_CDNS_756917543334 $T=64670 37880 0 0 $X=64530 $Y=37430
X203 8 VIA1_C_CDNS_756917543334 $T=64670 54100 0 0 $X=64530 $Y=53650
X204 11 VIA1_C_CDNS_756917543334 $T=64670 73000 0 0 $X=64530 $Y=72550
X205 11 VIA1_C_CDNS_756917543334 $T=65370 17120 0 0 $X=65230 $Y=16670
X206 11 VIA1_C_CDNS_756917543334 $T=65370 24340 0 0 $X=65230 $Y=23890
X207 11 VIA1_C_CDNS_756917543334 $T=65370 40560 0 0 $X=65230 $Y=40110
X208 11 VIA1_C_CDNS_756917543334 $T=65370 56780 0 0 $X=65230 $Y=56330
X209 11 VIA1_C_CDNS_756917543334 $T=65370 73000 0 0 $X=65230 $Y=72550
X210 11 VIA1_C_CDNS_756917543334 $T=66640 24340 0 0 $X=66500 $Y=23890
X211 5 VIA1_C_CDNS_756917543334 $T=66640 36540 0 0 $X=66500 $Y=36090
X212 5 VIA1_C_CDNS_756917543334 $T=66640 52760 0 0 $X=66500 $Y=52310
X213 5 VIA1_C_CDNS_756917543334 $T=66640 68980 0 0 $X=66500 $Y=68530
X214 11 VIA1_C_CDNS_756917543334 $T=67910 17120 0 0 $X=67770 $Y=16670
X215 8 VIA1_C_CDNS_756917543334 $T=67910 21660 0 0 $X=67770 $Y=21210
X216 8 VIA1_C_CDNS_756917543334 $T=67910 37880 0 0 $X=67770 $Y=37430
X217 8 VIA1_C_CDNS_756917543334 $T=67910 54100 0 0 $X=67770 $Y=53650
X218 11 VIA1_C_CDNS_756917543334 $T=67910 73000 0 0 $X=67770 $Y=72550
X219 11 VIA1_C_CDNS_756917543334 $T=68610 17120 0 0 $X=68470 $Y=16670
X220 11 VIA1_C_CDNS_756917543334 $T=68610 24340 0 0 $X=68470 $Y=23890
X221 11 VIA1_C_CDNS_756917543334 $T=68610 40560 0 0 $X=68470 $Y=40110
X222 11 VIA1_C_CDNS_756917543334 $T=68610 56780 0 0 $X=68470 $Y=56330
X223 11 VIA1_C_CDNS_756917543334 $T=68610 73000 0 0 $X=68470 $Y=72550
X224 11 VIA1_C_CDNS_756917543334 $T=69880 24340 0 0 $X=69740 $Y=23890
X225 5 VIA1_C_CDNS_756917543334 $T=69880 36540 0 0 $X=69740 $Y=36090
X226 5 VIA1_C_CDNS_756917543334 $T=69880 52760 0 0 $X=69740 $Y=52310
X227 5 VIA1_C_CDNS_756917543334 $T=69880 68980 0 0 $X=69740 $Y=68530
X228 11 VIA1_C_CDNS_756917543334 $T=71150 17120 0 0 $X=71010 $Y=16670
X229 8 VIA1_C_CDNS_756917543334 $T=71150 21660 0 0 $X=71010 $Y=21210
X230 8 VIA1_C_CDNS_756917543334 $T=71150 37880 0 0 $X=71010 $Y=37430
X231 8 VIA1_C_CDNS_756917543334 $T=71150 54100 0 0 $X=71010 $Y=53650
X232 11 VIA1_C_CDNS_756917543334 $T=71150 73000 0 0 $X=71010 $Y=72550
X233 11 VIA1_C_CDNS_756917543334 $T=71850 17120 0 0 $X=71710 $Y=16670
X234 11 VIA1_C_CDNS_756917543334 $T=71850 24340 0 0 $X=71710 $Y=23890
X235 11 VIA1_C_CDNS_756917543334 $T=71850 40560 0 0 $X=71710 $Y=40110
X236 11 VIA1_C_CDNS_756917543334 $T=71850 56780 0 0 $X=71710 $Y=56330
X237 11 VIA1_C_CDNS_756917543334 $T=71850 73000 0 0 $X=71710 $Y=72550
X238 11 VIA1_C_CDNS_756917543334 $T=73120 24340 0 0 $X=72980 $Y=23890
X239 5 VIA1_C_CDNS_756917543334 $T=73120 36540 0 0 $X=72980 $Y=36090
X240 5 VIA1_C_CDNS_756917543334 $T=73120 52760 0 0 $X=72980 $Y=52310
X241 5 VIA1_C_CDNS_756917543334 $T=73120 68980 0 0 $X=72980 $Y=68530
X242 11 VIA1_C_CDNS_756917543334 $T=74390 17120 0 0 $X=74250 $Y=16670
X243 8 VIA1_C_CDNS_756917543334 $T=74390 21660 0 0 $X=74250 $Y=21210
X244 8 VIA1_C_CDNS_756917543334 $T=74390 37880 0 0 $X=74250 $Y=37430
X245 8 VIA1_C_CDNS_756917543334 $T=74390 54100 0 0 $X=74250 $Y=53650
X246 11 VIA1_C_CDNS_756917543334 $T=74390 73000 0 0 $X=74250 $Y=72550
X247 11 VIA1_C_CDNS_756917543334 $T=75090 24340 0 0 $X=74950 $Y=23890
X248 11 VIA1_C_CDNS_756917543334 $T=75090 40560 0 0 $X=74950 $Y=40110
X249 11 VIA1_C_CDNS_756917543334 $T=75090 56780 0 0 $X=74950 $Y=56330
X250 11 VIA1_C_CDNS_756917543334 $T=75090 73000 0 0 $X=74950 $Y=72550
X251 11 VIA1_C_CDNS_756917543334 $T=76360 17120 0 0 $X=76220 $Y=16670
X252 5 VIA1_C_CDNS_756917543334 $T=76360 36540 0 0 $X=76220 $Y=36090
X253 5 VIA1_C_CDNS_756917543334 $T=76360 52760 0 0 $X=76220 $Y=52310
X254 5 VIA1_C_CDNS_756917543334 $T=76360 68980 0 0 $X=76220 $Y=68530
X255 7 VIA1_C_CDNS_756917543334 $T=77630 23000 0 0 $X=77490 $Y=22550
X256 5 VIA1_C_CDNS_756917543334 $T=77630 36540 0 0 $X=77490 $Y=36090
X257 7 VIA1_C_CDNS_756917543334 $T=77630 55440 0 0 $X=77490 $Y=54990
X258 11 VIA1_C_CDNS_756917543334 $T=77630 73000 0 0 $X=77490 $Y=72550
X259 11 VIA1_C_CDNS_756917543334 $T=78200 17120 0 0 $X=78060 $Y=16670
X260 11 VIA1_C_CDNS_756917543334 $T=78330 24340 0 0 $X=78190 $Y=23890
X261 11 VIA1_C_CDNS_756917543334 $T=78330 40560 0 0 $X=78190 $Y=40110
X262 11 VIA1_C_CDNS_756917543334 $T=78330 56780 0 0 $X=78190 $Y=56330
X263 11 VIA1_C_CDNS_756917543334 $T=78330 73000 0 0 $X=78190 $Y=72550
X264 11 VIA1_C_CDNS_756917543334 $T=79600 24340 0 0 $X=79460 $Y=23890
X265 5 VIA1_C_CDNS_756917543334 $T=79600 36540 0 0 $X=79460 $Y=36090
X266 5 VIA1_C_CDNS_756917543334 $T=79600 52760 0 0 $X=79460 $Y=52310
X267 5 VIA1_C_CDNS_756917543334 $T=79600 68980 0 0 $X=79460 $Y=68530
X268 11 VIA1_C_CDNS_756917543334 $T=80870 17120 0 0 $X=80730 $Y=16670
X269 7 VIA1_C_CDNS_756917543334 $T=80870 23000 0 0 $X=80730 $Y=22550
X270 5 VIA1_C_CDNS_756917543334 $T=80870 36540 0 0 $X=80730 $Y=36090
X271 7 VIA1_C_CDNS_756917543334 $T=80870 55440 0 0 $X=80730 $Y=54990
X272 11 VIA1_C_CDNS_756917543334 $T=80870 73000 0 0 $X=80730 $Y=72550
X273 11 VIA1_C_CDNS_756917543334 $T=81570 17120 0 0 $X=81430 $Y=16670
X274 11 VIA1_C_CDNS_756917543334 $T=81570 24340 0 0 $X=81430 $Y=23890
X275 11 VIA1_C_CDNS_756917543334 $T=81570 40560 0 0 $X=81430 $Y=40110
X276 11 VIA1_C_CDNS_756917543334 $T=81570 56780 0 0 $X=81430 $Y=56330
X277 11 VIA1_C_CDNS_756917543334 $T=81570 73000 0 0 $X=81430 $Y=72550
X278 11 VIA1_C_CDNS_756917543334 $T=82840 24340 0 0 $X=82700 $Y=23890
X279 5 VIA1_C_CDNS_756917543334 $T=82840 36540 0 0 $X=82700 $Y=36090
X280 5 VIA1_C_CDNS_756917543334 $T=82840 52760 0 0 $X=82700 $Y=52310
X281 5 VIA1_C_CDNS_756917543334 $T=82840 68980 0 0 $X=82700 $Y=68530
X282 11 VIA1_C_CDNS_756917543334 $T=84110 17120 0 0 $X=83970 $Y=16670
X283 8 VIA1_C_CDNS_756917543334 $T=84110 21660 0 0 $X=83970 $Y=21210
X284 8 VIA1_C_CDNS_756917543334 $T=84110 37880 0 0 $X=83970 $Y=37430
X285 8 VIA1_C_CDNS_756917543334 $T=84110 54100 0 0 $X=83970 $Y=53650
X286 11 VIA1_C_CDNS_756917543334 $T=84110 73000 0 0 $X=83970 $Y=72550
X287 11 VIA1_C_CDNS_756917543334 $T=84810 17120 0 0 $X=84670 $Y=16670
X288 11 VIA1_C_CDNS_756917543334 $T=84810 24340 0 0 $X=84670 $Y=23890
X289 11 VIA1_C_CDNS_756917543334 $T=84810 40560 0 0 $X=84670 $Y=40110
X290 11 VIA1_C_CDNS_756917543334 $T=84810 56780 0 0 $X=84670 $Y=56330
X291 11 VIA1_C_CDNS_756917543334 $T=84810 73000 0 0 $X=84670 $Y=72550
X292 11 VIA1_C_CDNS_756917543334 $T=86080 24340 0 0 $X=85940 $Y=23890
X293 5 VIA1_C_CDNS_756917543334 $T=86080 36540 0 0 $X=85940 $Y=36090
X294 5 VIA1_C_CDNS_756917543334 $T=86080 52760 0 0 $X=85940 $Y=52310
X295 5 VIA1_C_CDNS_756917543334 $T=86080 68980 0 0 $X=85940 $Y=68530
X296 11 VIA1_C_CDNS_756917543334 $T=87350 17120 0 0 $X=87210 $Y=16670
X297 8 VIA1_C_CDNS_756917543334 $T=87350 21660 0 0 $X=87210 $Y=21210
X298 8 VIA1_C_CDNS_756917543334 $T=87350 37880 0 0 $X=87210 $Y=37430
X299 8 VIA1_C_CDNS_756917543334 $T=87350 54100 0 0 $X=87210 $Y=53650
X300 11 VIA1_C_CDNS_756917543334 $T=87350 73000 0 0 $X=87210 $Y=72550
X301 11 VIA1_C_CDNS_756917543334 $T=88050 17120 0 0 $X=87910 $Y=16670
X302 11 VIA1_C_CDNS_756917543334 $T=88050 24340 0 0 $X=87910 $Y=23890
X303 11 VIA1_C_CDNS_756917543334 $T=88050 40560 0 0 $X=87910 $Y=40110
X304 11 VIA1_C_CDNS_756917543334 $T=88050 56780 0 0 $X=87910 $Y=56330
X305 11 VIA1_C_CDNS_756917543334 $T=88050 73000 0 0 $X=87910 $Y=72550
X306 11 VIA1_C_CDNS_756917543334 $T=89320 24340 0 0 $X=89180 $Y=23890
X307 5 VIA1_C_CDNS_756917543334 $T=89320 36540 0 0 $X=89180 $Y=36090
X308 5 VIA1_C_CDNS_756917543334 $T=89320 52760 0 0 $X=89180 $Y=52310
X309 5 VIA1_C_CDNS_756917543334 $T=89320 68980 0 0 $X=89180 $Y=68530
X310 11 VIA1_C_CDNS_756917543334 $T=90590 17120 0 0 $X=90450 $Y=16670
X311 8 VIA1_C_CDNS_756917543334 $T=90590 21660 0 0 $X=90450 $Y=21210
X312 8 VIA1_C_CDNS_756917543334 $T=90590 37880 0 0 $X=90450 $Y=37430
X313 8 VIA1_C_CDNS_756917543334 $T=90590 54100 0 0 $X=90450 $Y=53650
X314 11 VIA1_C_CDNS_756917543334 $T=90590 73000 0 0 $X=90450 $Y=72550
X315 11 VIA1_C_CDNS_756917543334 $T=91290 17120 0 0 $X=91150 $Y=16670
X316 11 VIA1_C_CDNS_756917543334 $T=91290 24340 0 0 $X=91150 $Y=23890
X317 11 VIA1_C_CDNS_756917543334 $T=91290 40560 0 0 $X=91150 $Y=40110
X318 11 VIA1_C_CDNS_756917543334 $T=91290 56780 0 0 $X=91150 $Y=56330
X319 11 VIA1_C_CDNS_756917543334 $T=91290 73000 0 0 $X=91150 $Y=72550
X320 11 VIA1_C_CDNS_756917543334 $T=92560 24340 0 0 $X=92420 $Y=23890
X321 5 VIA1_C_CDNS_756917543334 $T=92560 36540 0 0 $X=92420 $Y=36090
X322 5 VIA1_C_CDNS_756917543334 $T=92560 52760 0 0 $X=92420 $Y=52310
X323 5 VIA1_C_CDNS_756917543334 $T=92560 68980 0 0 $X=92420 $Y=68530
X324 11 VIA1_C_CDNS_756917543334 $T=93830 17120 0 0 $X=93690 $Y=16670
X325 8 VIA1_C_CDNS_756917543334 $T=93830 21660 0 0 $X=93690 $Y=21210
X326 8 VIA1_C_CDNS_756917543334 $T=93830 37880 0 0 $X=93690 $Y=37430
X327 8 VIA1_C_CDNS_756917543334 $T=93830 54100 0 0 $X=93690 $Y=53650
X328 11 VIA1_C_CDNS_756917543334 $T=93830 73000 0 0 $X=93690 $Y=72550
X329 11 VIA1_C_CDNS_756917543334 $T=94530 17120 0 0 $X=94390 $Y=16670
X330 11 VIA1_C_CDNS_756917543334 $T=94530 24340 0 0 $X=94390 $Y=23890
X331 11 VIA1_C_CDNS_756917543334 $T=94530 40560 0 0 $X=94390 $Y=40110
X332 11 VIA1_C_CDNS_756917543334 $T=94530 56780 0 0 $X=94390 $Y=56330
X333 11 VIA1_C_CDNS_756917543334 $T=94530 73000 0 0 $X=94390 $Y=72550
X334 11 VIA1_C_CDNS_756917543334 $T=95800 24340 0 0 $X=95660 $Y=23890
X335 5 VIA1_C_CDNS_756917543334 $T=95800 36540 0 0 $X=95660 $Y=36090
X336 5 VIA1_C_CDNS_756917543334 $T=95800 52760 0 0 $X=95660 $Y=52310
X337 5 VIA1_C_CDNS_756917543334 $T=95800 68980 0 0 $X=95660 $Y=68530
X338 11 VIA1_C_CDNS_756917543334 $T=97070 17120 0 0 $X=96930 $Y=16670
X339 8 VIA1_C_CDNS_756917543334 $T=97070 21660 0 0 $X=96930 $Y=21210
X340 8 VIA1_C_CDNS_756917543334 $T=97070 37880 0 0 $X=96930 $Y=37430
X341 8 VIA1_C_CDNS_756917543334 $T=97070 54100 0 0 $X=96930 $Y=53650
X342 11 VIA1_C_CDNS_756917543334 $T=97070 73000 0 0 $X=96930 $Y=72550
X343 11 VIA1_C_CDNS_756917543334 $T=97770 17120 0 0 $X=97630 $Y=16670
X344 11 VIA1_C_CDNS_756917543334 $T=97770 24340 0 0 $X=97630 $Y=23890
X345 11 VIA1_C_CDNS_756917543334 $T=97770 40560 0 0 $X=97630 $Y=40110
X346 11 VIA1_C_CDNS_756917543334 $T=97770 56780 0 0 $X=97630 $Y=56330
X347 11 VIA1_C_CDNS_756917543334 $T=97770 73000 0 0 $X=97630 $Y=72550
X348 11 VIA1_C_CDNS_756917543334 $T=99040 24340 0 0 $X=98900 $Y=23890
X349 11 VIA1_C_CDNS_756917543334 $T=99040 40560 0 0 $X=98900 $Y=40110
X350 11 VIA1_C_CDNS_756917543334 $T=99040 56780 0 0 $X=98900 $Y=56330
X351 11 VIA1_C_CDNS_756917543334 $T=99040 73000 0 0 $X=98900 $Y=72550
X352 11 VIA1_C_CDNS_756917543334 $T=100310 17120 0 0 $X=100170 $Y=16670
X353 11 VIA1_C_CDNS_756917543334 $T=100310 24340 0 0 $X=100170 $Y=23890
X354 11 VIA1_C_CDNS_756917543334 $T=100310 40560 0 0 $X=100170 $Y=40110
X355 11 VIA1_C_CDNS_756917543334 $T=100310 56780 0 0 $X=100170 $Y=56330
X356 11 VIA1_C_CDNS_756917543334 $T=100310 73000 0 0 $X=100170 $Y=72550
X357 5 VIA2_C_CDNS_756917543336 $T=50410 13100 0 0 $X=49700 $Y=12700
X358 5 VIA2_C_CDNS_756917543336 $T=50410 20320 0 0 $X=49700 $Y=19920
X359 5 VIA2_C_CDNS_756917543336 $T=50410 36540 0 0 $X=49700 $Y=36140
X360 5 VIA2_C_CDNS_756917543336 $T=50410 52760 0 0 $X=49700 $Y=52360
X361 5 VIA2_C_CDNS_756917543336 $T=50410 68980 0 0 $X=49700 $Y=68580
X362 7 VIA2_C_CDNS_756917543336 $T=52250 15780 0 0 $X=51540 $Y=15380
X363 7 VIA2_C_CDNS_756917543336 $T=52250 23000 0 0 $X=51540 $Y=22600
X364 7 VIA2_C_CDNS_756917543336 $T=52250 39220 0 0 $X=51540 $Y=38820
X365 7 VIA2_C_CDNS_756917543336 $T=52250 55440 0 0 $X=51540 $Y=55040
X366 7 VIA2_C_CDNS_756917543336 $T=52250 71660 0 0 $X=51540 $Y=71260
X367 11 VIA2_C_CDNS_756917543336 $T=54090 17120 0 0 $X=53380 $Y=16720
X368 11 VIA2_C_CDNS_756917543336 $T=54090 24340 0 0 $X=53380 $Y=23940
X369 11 VIA2_C_CDNS_756917543336 $T=54090 40560 0 0 $X=53380 $Y=40160
X370 11 VIA2_C_CDNS_756917543336 $T=54090 56780 0 0 $X=53380 $Y=56380
X371 11 VIA2_C_CDNS_756917543336 $T=54090 73000 0 0 $X=53380 $Y=72600
X372 11 VIA2_C_CDNS_756917543336 $T=101870 17120 0 0 $X=101160 $Y=16720
X373 11 VIA2_C_CDNS_756917543336 $T=101870 24340 0 0 $X=101160 $Y=23940
X374 11 VIA2_C_CDNS_756917543336 $T=101870 40560 0 0 $X=101160 $Y=40160
X375 11 VIA2_C_CDNS_756917543336 $T=101870 56780 0 0 $X=101160 $Y=56380
X376 11 VIA2_C_CDNS_756917543336 $T=101870 73000 0 0 $X=101160 $Y=72600
X377 8 VIA2_C_CDNS_756917543336 $T=103710 14440 0 0 $X=103000 $Y=14040
X378 8 VIA2_C_CDNS_756917543336 $T=103710 21660 0 0 $X=103000 $Y=21260
X379 8 VIA2_C_CDNS_756917543336 $T=103710 37880 0 0 $X=103000 $Y=37480
X380 8 VIA2_C_CDNS_756917543336 $T=103710 54100 0 0 $X=103000 $Y=53700
X381 8 VIA2_C_CDNS_756917543336 $T=103710 70320 0 0 $X=103000 $Y=69920
X382 6 VIA1_C_CDNS_756917543338 $T=7520 29745 0 0 $X=6510 $Y=28995
X383 1 VIA1_C_CDNS_756917543338 $T=61555 108745 0 0 $X=60545 $Y=107995
X384 1 VIA1_C_CDNS_756917543338 $T=68285 108255 0 0 $X=67275 $Y=107505
X385 6 VIA1_C_CDNS_756917543339 $T=25375 26765 0 0 $X=24365 $Y=26275
X386 2 VIA1_C_CDNS_756917543339 $T=50500 95625 0 0 $X=49490 $Y=95135
X387 2 VIA1_C_CDNS_756917543339 $T=53560 100075 0 0 $X=52550 $Y=99585
X388 12 VIA1_C_CDNS_756917543339 $T=70840 95455 0 0 $X=69830 $Y=94965
X389 7 VIA2_C_CDNS_7569175433317 $T=52250 29260 0 0 $X=51500 $Y=28510
X390 8 VIA2_C_CDNS_7569175433317 $T=53535 106615 0 0 $X=52785 $Y=105865
X391 2 12 1 11 rpp1k1_3_CDNS_756917543330 $T=71840 92685 1 270 $X=49280 $Y=80495
X392 7 6 4 11 nel_CDNS_756917543331 $T=31115 23480 1 0 $X=30375 $Y=17910
X393 5 6 11 nel_CDNS_756917543332 $T=18470 23480 1 0 $X=17730 $Y=17910
X394 1 2 8 11 pel_CDNS_756917543334 $T=57470 103255 0 180 $X=48780 $Y=100185
X395 11 11 11 11 nel_CDNS_756917543335 $T=12080 38620 0 0 $X=11340 $Y=38270
X396 11 11 11 11 nel_CDNS_756917543335 $T=12080 61580 1 0 $X=11340 $Y=51010
X397 4 9 3 11 nel_CDNS_756917543335 $T=14320 38620 0 0 $X=13580 $Y=38270
X398 4 10 2 11 nel_CDNS_756917543335 $T=14320 61580 1 0 $X=13580 $Y=51010
X399 4 10 2 11 nel_CDNS_756917543335 $T=16560 38620 0 0 $X=15820 $Y=38270
X400 4 9 3 11 nel_CDNS_756917543335 $T=16560 61580 1 0 $X=15820 $Y=51010
X401 4 9 3 11 nel_CDNS_756917543335 $T=18800 38620 0 0 $X=18060 $Y=38270
X402 4 10 2 11 nel_CDNS_756917543335 $T=18800 61580 1 0 $X=18060 $Y=51010
X403 4 10 2 11 nel_CDNS_756917543335 $T=21040 38620 0 0 $X=20300 $Y=38270
X404 4 9 3 11 nel_CDNS_756917543335 $T=21040 61580 1 0 $X=20300 $Y=51010
X405 4 9 3 11 nel_CDNS_756917543335 $T=23280 38620 0 0 $X=22540 $Y=38270
X406 4 10 2 11 nel_CDNS_756917543335 $T=23280 61580 1 0 $X=22540 $Y=51010
X407 4 10 2 11 nel_CDNS_756917543335 $T=25520 38620 0 0 $X=24780 $Y=38270
X408 4 9 3 11 nel_CDNS_756917543335 $T=25520 61580 1 0 $X=24780 $Y=51010
X409 4 9 3 11 nel_CDNS_756917543335 $T=27760 38620 0 0 $X=27020 $Y=38270
X410 4 10 2 11 nel_CDNS_756917543335 $T=27760 61580 1 0 $X=27020 $Y=51010
X411 4 10 2 11 nel_CDNS_756917543335 $T=30000 38620 0 0 $X=29260 $Y=38270
X412 4 9 3 11 nel_CDNS_756917543335 $T=30000 61580 1 0 $X=29260 $Y=51010
X413 4 9 3 11 nel_CDNS_756917543335 $T=32240 38620 0 0 $X=31500 $Y=38270
X414 4 10 2 11 nel_CDNS_756917543335 $T=32240 61580 1 0 $X=31500 $Y=51010
X415 4 10 2 11 nel_CDNS_756917543335 $T=34480 38620 0 0 $X=33740 $Y=38270
X416 4 9 3 11 nel_CDNS_756917543335 $T=34480 61580 1 0 $X=33740 $Y=51010
X417 11 11 11 11 nel_CDNS_756917543335 $T=36720 38620 0 0 $X=35980 $Y=38270
X418 11 11 11 11 nel_CDNS_756917543335 $T=36720 61580 1 0 $X=35980 $Y=51010
X419 1 1 1 11 pel_CDNS_756917543336 $T=8410 79155 0 0 $X=7500 $Y=78725
X420 1 1 1 11 pel_CDNS_756917543336 $T=8410 101415 1 0 $X=7500 $Y=90845
X421 1 3 2 11 pel_CDNS_756917543336 $T=11650 79155 0 0 $X=10740 $Y=78725
X422 1 3 3 11 pel_CDNS_756917543336 $T=11650 101415 1 0 $X=10740 $Y=90845
X423 1 3 3 11 pel_CDNS_756917543336 $T=14890 79155 0 0 $X=13980 $Y=78725
X424 1 3 2 11 pel_CDNS_756917543336 $T=14890 101415 1 0 $X=13980 $Y=90845
X425 1 3 2 11 pel_CDNS_756917543336 $T=18130 79155 0 0 $X=17220 $Y=78725
X426 1 3 3 11 pel_CDNS_756917543336 $T=18130 101415 1 0 $X=17220 $Y=90845
X427 1 3 3 11 pel_CDNS_756917543336 $T=21370 79155 0 0 $X=20460 $Y=78725
X428 1 3 2 11 pel_CDNS_756917543336 $T=21370 101415 1 0 $X=20460 $Y=90845
X429 1 3 3 11 pel_CDNS_756917543336 $T=24610 79155 0 0 $X=23700 $Y=78725
X430 1 3 2 11 pel_CDNS_756917543336 $T=24610 101415 1 0 $X=23700 $Y=90845
X431 1 3 2 11 pel_CDNS_756917543336 $T=27850 79155 0 0 $X=26940 $Y=78725
X432 1 3 3 11 pel_CDNS_756917543336 $T=27850 101415 1 0 $X=26940 $Y=90845
X433 1 3 3 11 pel_CDNS_756917543336 $T=31090 79155 0 0 $X=30180 $Y=78725
X434 1 3 2 11 pel_CDNS_756917543336 $T=31090 101415 1 0 $X=30180 $Y=90845
X435 1 3 2 11 pel_CDNS_756917543336 $T=34330 79155 0 0 $X=33420 $Y=78725
X436 1 3 3 11 pel_CDNS_756917543336 $T=34330 101415 1 0 $X=33420 $Y=90845
X437 1 1 1 11 pel_CDNS_756917543336 $T=37570 79155 0 0 $X=36660 $Y=78725
X438 1 1 1 11 pel_CDNS_756917543336 $T=37570 101415 1 0 $X=36660 $Y=90845
X439 11 1 mosvc_CDNS_756917543339 $T=63350 99890 0 0 $X=62610 $Y=99460
X440 11 6 mosvc_CDNS_7569175433310 $T=2695 11965 0 0 $X=1955 $Y=11535
X441 11 MASCO__A1 $T=55180 17760 0 0 $X=55180 $Y=17760
X442 11 MASCO__A1 $T=55180 73640 0 0 $X=55180 $Y=73640
X443 11 MASCO__A1 $T=61660 17760 0 0 $X=61660 $Y=17760
X444 11 MASCO__A1 $T=61660 73640 0 0 $X=61660 $Y=73640
X445 11 MASCO__A1 $T=68140 17760 0 0 $X=68140 $Y=17760
X446 11 MASCO__A1 $T=68140 73640 0 0 $X=68140 $Y=73640
X447 11 MASCO__A1 $T=74620 17760 0 0 $X=74620 $Y=17760
X448 11 MASCO__A1 $T=74620 73640 0 0 $X=74620 $Y=73640
X449 11 MASCO__A1 $T=81100 17760 0 0 $X=81100 $Y=17760
X450 11 MASCO__A1 $T=81100 73640 0 0 $X=81100 $Y=73640
X451 11 MASCO__A1 $T=87580 17760 0 0 $X=87580 $Y=17760
X452 11 MASCO__A1 $T=87580 73640 0 0 $X=87580 $Y=73640
X453 11 MASCO__A1 $T=94060 17760 0 0 $X=94060 $Y=17760
X454 11 MASCO__A1 $T=94060 73640 0 0 $X=94060 $Y=73640
X455 11 5 8 11 11 MASCO__A2 $T=94060 24980 0 0 $X=94060 $Y=24980
X456 11 5 8 11 11 MASCO__A2 $T=94060 41200 0 0 $X=94060 $Y=41200
X457 11 5 8 11 11 MASCO__A2 $T=94060 57420 0 0 $X=94060 $Y=57420
X458 11 11 11 5 8 8 MASCO__A3 $T=55180 24980 0 0 $X=55180 $Y=24980
X459 11 11 11 5 8 8 MASCO__A3 $T=55180 41200 0 0 $X=55180 $Y=41200
X460 11 11 11 5 8 8 MASCO__A3 $T=55180 57420 0 0 $X=55180 $Y=57420
X461 11 5 8 5 8 7 MASCO__A3 $T=68140 24980 0 0 $X=68140 $Y=24980
X462 11 5 8 5 8 5 MASCO__A3 $T=68140 41200 0 0 $X=68140 $Y=41200
X463 11 5 8 5 8 7 MASCO__A3 $T=68140 57420 0 0 $X=68140 $Y=57420
X464 11 5 8 5 8 8 MASCO__A3 $T=81100 24980 0 0 $X=81100 $Y=24980
X465 11 5 8 5 8 8 MASCO__A3 $T=81100 41200 0 0 $X=81100 $Y=41200
X466 11 5 8 5 8 8 MASCO__A3 $T=81100 57420 0 0 $X=81100 $Y=57420
D0 11 1 p_dnw AREA=1.63313e-09 PJ=0.00016212 perimeter=0.00016212 $X=2180 $Y=71565 $dt=3
D1 11 1 p_dnw AREA=1.34725e-10 PJ=4.668e-05 perimeter=4.668e-05 $X=47140 $Y=98545 $dt=3
D2 11 1 p_dnw AREA=4.85498e-10 PJ=8.938e-05 perimeter=8.938e-05 $X=47640 $Y=78855 $dt=3
D3 11 1 p_dnw AREA=1.00372e-09 PJ=0.00012712 perimeter=0.00012712 $X=75350 $Y=79725 $dt=3
C4 12 8 area=7.5e-10 perimeter=0.00011 $[cmm5t] $X=77490 $Y=81865 $dt=5
.ends opamp1
